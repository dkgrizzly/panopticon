`timescale 1ns / 1ps
`default_nettype none
// Using 1 BRAM16_S1_S1
module bg0_map (
    input wire clka,
    input wire wea,
    input wire [13:0] addra,
    input wire dina,
    input wire clkb,
    input wire [13:0] addrb,
    output wire doutb
);

RAMB16_S1_S1 BRAM_BGMAP_0  (
  .CLKA(clka),
  .ENA(1'b1),
  .WEA(wea),
  .ADDRA(addra),
  .SSRA(1'b0),
  .DIA(dina),

  .CLKB(clkb),
  .ENB(1'b1),
  .WEB(1'b0),
  .ADDRB(addrb),
  .SSRB(1'b0),
  .DOB(doutb)
  );

defparam BRAM_BGMAP_0.INIT_00 = 256'h0050502751530107005050275457010700505077545701070000000000000000;
defparam BRAM_BGMAP_0.INIT_01 = 256'h0070101315130503005050355557050700207057517301070020202721730107;
defparam BRAM_BGMAP_0.INIT_02 = 256'h0020202225750505001010371171010100202025257705050070407315730503;
defparam BRAM_BGMAP_0.INIT_03 = 256'h0070202724770107007050575477010700503077517101070010103111730107;
defparam BRAM_BGMAP_0.INIT_04 = 256'h0070406345750503007010734575050300702023352505030070101315150503;
defparam BRAM_BGMAP_0.INIT_05 = 256'h0030503751330107002020775457010700505035555505070040407355550503;
defparam BRAM_BGMAP_0.INIT_06 = 256'h0070101711730107001800180C66663C00505057715301070050505751710107;
defparam BRAM_BGMAP_0.INIT_07 = 256'h0070407715750505007040751377050700704077157501070070407111730107;
defparam BRAM_BGMAP_0.INIT_08 = 256'h0036367F367F3636000000000066666600180018181818180000000000000000;
defparam BRAM_BGMAP_0.INIT_09 = 256'h00000000000C1818006E333B6E1C361C0063660C1833630000183E603C067C18;
defparam BRAM_BGMAP_0.INIT_0A = 256'h000018187E1818000000663CFF3C6600000C18303030180C0030180C0C0C1830;
defparam BRAM_BGMAP_0.INIT_0B = 256'h0003060C183060C00018180000000000000000007E0000000C18180000000000;
defparam BRAM_BGMAP_0.INIT_0C = 256'h003C66603860663C007E060C1830663C007E181818181C18003C66666E76663C;
defparam BRAM_BGMAP_0.INIT_0D = 256'h001818183060607E003C66663E060C38003C6660603E067E0030307F33363C38;
defparam BRAM_BGMAP_0.INIT_0E = 256'h0C181800001818000018180000181800001C30607C66663C003C66663C66663C;
defparam BRAM_BGMAP_0.INIT_0F = 256'h001800183060663C00060C1830180C060000007E007E00000030180C060C1830;
defparam BRAM_BGMAP_0.INIT_10 = 256'h003C66060606663C003E66663E66663E0066667E66663C18003E037B7B7B633E;
defparam BRAM_BGMAP_0.INIT_11 = 256'h007C66667606663C000606063E06067E007E06063E06067E001E36666666361E;
defparam BRAM_BGMAP_0.INIT_12 = 256'h0063331B0F1B3363003C666060606060007E18181818187E006666667E666666;
defparam BRAM_BGMAP_0.INIT_13 = 256'h003C66666666663C006363737B6F6763006363636B7F7763007E060606060606;
defparam BRAM_BGMAP_0.INIT_14 = 256'h003C66603C06663C006666363E66663E006C36666666663C000606063E66663E;
defparam BRAM_BGMAP_0.INIT_15 = 256'h0063777F6B63636300183C6666666666003C666666666666001818181818187E;
defparam BRAM_BGMAP_0.INIT_16 = 256'h003C0C0C0C0C0C3C007E060C1830607E00181818183C66C300C3663C183C66C3;
defparam BRAM_BGMAP_0.INIT_17 = 256'hFF000000000000000000000063361C08003C30303030303C00C06030180C0603;
defparam BRAM_BGMAP_0.INIT_18 = 256'h003C0606063C0000003E6666663E0606007C667C603C00000000000000603018;
defparam BRAM_BGMAP_0.INIT_19 = 256'h3E607C66667C0000000C0C0C0C3E0C38003C067E663C0000007C6666667C6060;
defparam BRAM_BGMAP_0.INIT_1A = 256'h0066361E366606061E3030303030003000781818181C001800666666663E0606;
defparam BRAM_BGMAP_0.INIT_1B = 256'h003C6666663C000000666666663E000000636B6B7F330000007818181818181C;
defparam BRAM_BGMAP_0.INIT_1C = 256'h003E603C067C000000060606663E000060607C66667C000006063E66663E0000;
defparam BRAM_BGMAP_0.INIT_1D = 256'h00363E6B6363000000183C6666660000007C66666666000000780C0C0C7E0C0C;
defparam BRAM_BGMAP_0.INIT_1E = 256'h007018180E181870007E0C18307E00003C607C66666600000063361C36630000;
defparam BRAM_BGMAP_0.INIT_1F = 256'h00202023257505030000000000003B6E000E18187018180E0018181818181818;
defparam BRAM_BGMAP_0.INIT_20 = 256'h0070407745770507007010774577050700702027352705070070505755770507;
defparam BRAM_BGMAP_0.INIT_21 = 256'h0070407711730107007040771477010700701015151505070050505752720207;
defparam BRAM_BGMAP_0.INIT_22 = 256'h0030505151370507007040721575050500705045454705050070407515770505;
defparam BRAM_BGMAP_0.INIT_23 = 256'h0070406744770107007010774477010700702025257305030070505151570507;
defparam BRAM_BGMAP_0.INIT_24 = 256'h0070103714770107007010714177050700702021312705070070101315750503;
defparam BRAM_BGMAP_0.INIT_25 = 256'h0010107751730107001010775477010700507075555707050070101711710107;
defparam BRAM_BGMAP_0.INIT_26 = 256'h0070407711710107005050775477050700704077547705070070507754770507;
defparam BRAM_BGMAP_0.INIT_27 = 256'h0010107555770507005050717157050700704077157505070020202724770107;
defparam BRAM_BGMAP_0.INIT_28 = 256'h003F66060F06361C00187E1B1B7E180000181818181800180000000000000000;
defparam BRAM_BGMAP_0.INIT_29 = 256'h3C603C66663C063C00181818001818180018183C183C66C3000000663C663C66;
defparam BRAM_BGMAP_0.INIT_2A = 256'h0000CC663366CC0000007E007C36363C7E81B98D8DB9817E0000000000000066;
defparam BRAM_BGMAP_0.INIT_2B = 256'h000000000000007E7E81A59DA59D817E000000003C0000000000000060607E00;
defparam BRAM_BGMAP_0.INIT_2C = 256'h0000001E3018301E0000001E060C180E007E0018187E181800000000003C663C;
defparam BRAM_BGMAP_0.INIT_2D = 256'h0000000018000000005858585C5E5E7C03063E666666000000000000000C1830;
defparam BRAM_BGMAP_0.INIT_2E = 256'h00003366CC66330000003E001C36361C0000000C0C0C0E0C1810000000000000;
defparam BRAM_BGMAP_0.INIT_2F = 256'h003C66060C18001840F3566F5C366403F03366CC7A32630240F3566C5A326302;
defparam BRAM_BGMAP_0.INIT_30 = 256'h00667E663C003B6E00667E663C0066180066667E663C00700066667E663C000E;
defparam BRAM_BGMAP_0.INIT_31 = 256'h183C66060606663C00F333337F3336FC00667E663C0018180066667E663C0066;
defparam BRAM_BGMAP_0.INIT_32 = 256'h007F031F037F0066007F030F7F006618007F031F037F0070007F031F037F000E;
defparam BRAM_BGMAP_0.INIT_33 = 256'h007E1818187E0066007E18187E006618007E1818187E0070007E1818187E000E;
defparam BRAM_BGMAP_0.INIT_34 = 256'h003E6363633E0070003E6363633E000E00637B6F63003B6E001E36666F66361E;
defparam BRAM_BGMAP_0.INIT_35 = 256'h000063361C366300003E6363633E0066003E63633E003B6E003E63633E006618;
defparam BRAM_BGMAP_0.INIT_36 = 256'h003E636363006618003E636363630070003E63636363000E003E666E7E76667C;
defparam BRAM_BGMAP_0.INIT_37 = 256'h003666663666663C0003033F633F03030018183C66660070003E636363630066;
defparam BRAM_BGMAP_0.INIT_38 = 256'h007E63667C003B6E007E63667C006618007C667C603C0070007C667C603C000E;
defparam BRAM_BGMAP_0.INIT_39 = 256'h183C0606063C000000EE1BFED87E0000007E63667C001818007C667C603C0066;
defparam BRAM_BGMAP_0.INIT_3A = 256'h003C067E663C0066003C067E3C006618003C067E663C0070003C067E663C000E;
defparam BRAM_BGMAP_0.INIT_3B = 256'h003C1818181C0066003C18181C006618003C1818181C0070003C1818181C000E;
defparam BRAM_BGMAP_0.INIT_3C = 256'h003C6666663C0070003C6666663C000E006666663E003B6E001E33333E307C30;
defparam BRAM_BGMAP_0.INIT_3D = 256'h001818007E001818003C6666663C0066003C66663C003B6E003C66663C006618;
defparam BRAM_BGMAP_0.INIT_3E = 256'h007C666666006618007C666666660070007C66666666000E013E676B733E4000;
defparam BRAM_BGMAP_0.INIT_3F = 256'h3C607C666666006606063E66663E06063C607C6666660070007C666666660066;
endmodule
