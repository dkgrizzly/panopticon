// Palette RAM 512x32 XRGB - Using 1 BRAM16_S36_S36
`timescale 1ns / 1ps
`default_nettype none
module palette_ram (
    input wire clka,
    input wire wea,
    input wire [8:0] addra,
    input wire [31:0] dina,
    input wire clkb,
    input wire [8:0] addrb,
    output wire [31:0] doutb
);

RAMB16_S36_S36 BRAM_PALMAP_0  (
  .CLKA(clka),
  .ENA(1'b1),
  .WEA(wea),
  .ADDRA(addra),
  .SSRA(1'b0),
  .DIA(dina),
  .DIPA(4'd0),

  .CLKB(clkb),
  .ENB(1'b1),
  .WEB(1'b0),
  .ADDRB(addrb),
  .SSRB(1'b0),
  .DOB(doutb)
  );

defparam BRAM_PALMAP_0.INIT_00 = 256'h0303030001010000010001000100000000010100000100000000010000000000;
defparam BRAM_PALMAP_0.INIT_01 = 256'hFFFFFF00FFFF0000FF00FF00FF00000000FFFF0000FF00000000FF0001010100;
defparam BRAM_PALMAP_0.INIT_02 = 256'hFAFA000000FA0000FF000000EB000000F5000000E1000000FA00000000000000;
defparam BRAM_PALMAP_0.INIT_03 = 256'hF5E10000E1E10000FAE1000000E10000FFFA0000EBFA0000F5FA0000E1FA0000;
defparam BRAM_PALMAP_0.INIT_04 = 256'hFFF50000EBF50000F5F50000E1F50000FAF5000000F50000FFE10000EBE10000;
defparam BRAM_PALMAP_0.INIT_05 = 256'hFAFF000000FF0000FFEB0000EBEB0000F5EB0000E1EB0000FAEB000000EB0000;
defparam BRAM_PALMAP_0.INIT_06 = 256'hF500FA00E100FA00FA00FA000000FA00FFFF0000EBFF0000F5FF0000E1FF0000;
defparam BRAM_PALMAP_0.INIT_07 = 256'hFFFAFA00EBFAFA00F5FAFA00E1FAFA00FAFAFA0000FAFA00FF00FA00EB00FA00;
defparam BRAM_PALMAP_0.INIT_08 = 256'hFAF5FA0000F5FA00FFE1FA00EBE1FA00F5E1FA00E1E1FA00FAE1FA0000E1FA00;
defparam BRAM_PALMAP_0.INIT_09 = 256'hF5EBFA00E1EBFA00FAEBFA0000EBFA00FFF5FA00EBF5FA00F5F5FA00E1F5FA00;
defparam BRAM_PALMAP_0.INIT_0A = 256'hFFFFFA00EBFFFA00F5FFFA00E1FFFA00FAFFFA0000FFFA00FFEBFA00EBEBFA00;
defparam BRAM_PALMAP_0.INIT_0B = 256'hFAFAE10000FAE100FF00E100EB00E100F500E100E100E100FA00E1000000E100;
defparam BRAM_PALMAP_0.INIT_0C = 256'hF5E1E100E1E1E100FAE1E10000E1E100FFFAE100EBFAE100F5FAE100E1FAE100;
defparam BRAM_PALMAP_0.INIT_0D = 256'hFFF5E100EBF5E100F5F5E100E1F5E100FAF5E10000F5E100FFE1E100EBE1E100;
defparam BRAM_PALMAP_0.INIT_0E = 256'hFAFFE10000FFE100FFEBE100EBEBE100F5EBE100E1EBE100FAEBE10000EBE100;
defparam BRAM_PALMAP_0.INIT_0F = 256'hF500F500E100F500FA00F5000000F500FFFFE100EBFFE100F5FFE100E1FFE100;
defparam BRAM_PALMAP_0.INIT_10 = 256'hFFFAF500EBFAF500F5FAF500E1FAF500FAFAF50000FAF500FF00F500EB00F500;
defparam BRAM_PALMAP_0.INIT_11 = 256'hFAF5F50000F5F500FFE1F500EBE1F500F5E1F500E1E1F500FAE1F50000E1F500;
defparam BRAM_PALMAP_0.INIT_12 = 256'hF5EBF500E1EBF500FAEBF50000EBF500FFF5F500EBF5F500F5F5F500E1F5F500;
defparam BRAM_PALMAP_0.INIT_13 = 256'hFFFFF500EBFFF500F5FFF500E1FFF500FAFFF50000FFF500FFEBF500EBEBF500;
defparam BRAM_PALMAP_0.INIT_14 = 256'hFAFAEB0000FAEB00FF00EB00EB00EB00F500EB00E100EB00FA00EB000000EB00;
defparam BRAM_PALMAP_0.INIT_15 = 256'hF5E1EB00E1E1EB00FAE1EB0000E1EB00FFFAEB00EBFAEB00F5FAEB00E1FAEB00;
defparam BRAM_PALMAP_0.INIT_16 = 256'hFFF5EB00EBF5EB00F5F5EB00E1F5EB00FAF5EB0000F5EB00FFE1EB00EBE1EB00;
defparam BRAM_PALMAP_0.INIT_17 = 256'hFAFFEB0000FFEB00FFEBEB00EBEBEB00F5EBEB00E1EBEB00FAEBEB0000EBEB00;
defparam BRAM_PALMAP_0.INIT_18 = 256'hF500FF00E100FF00FA00FF000000FF00FFFFEB00EBFFEB00F5FFEB00E1FFEB00;
defparam BRAM_PALMAP_0.INIT_19 = 256'hFFFAFF00EBFAFF00F5FAFF00E1FAFF00FAFAFF0000FAFF00FF00FF00EB00FF00;
defparam BRAM_PALMAP_0.INIT_1A = 256'hFAF5FF0000F5FF00FFE1FF00EBE1FF00F5E1FF00E1E1FF00FAE1FF0000E1FF00;
defparam BRAM_PALMAP_0.INIT_1B = 256'hF5EBFF00E1EBFF00FAEBFF0000EBFF00FFF5FF00EBF5FF00F5F5FF00E1F5FF00;
defparam BRAM_PALMAP_0.INIT_1C = 256'hFFFFFF00EBFFFF00F5FFFF00E1FFFF00FAFFFF0000FFFF00FFEBFF00EBEBFF00;
defparam BRAM_PALMAP_0.INIT_1D = 256'h72727200222222005C5C5C000C0C0C0064646400383838004848480010101000;
defparam BRAM_PALMAP_0.INIT_1E = 256'h797979002929290051515100010101006E6E6E0036363600464646001A1A1A00;
defparam BRAM_PALMAP_0.INIT_1F = 256'h77777700272727005B5B5B000B0B0B00636363003D3D3D004D4D4D0015151500;

endmodule
