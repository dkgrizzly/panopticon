`timescale 1ns / 1ps
`default_nettype none
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Wenting Zhang
// 
// Create Date:    15:28:43 02/07/2018 
// Design Name: 
// Module Name:    vga_mixer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vga_mixer(
    input wire vga_clk,
    input wire vga_rst,
    
    // CPU Bus Interface
    input wire cpu_clk,
    input wire vga_reg_wea,
    input wire vga_pal_wea,
    input wire vga_cop_wea,
    input wire vga_oam_wea,
    input wire vga_spr_wea,
    input wire vga_bt0_wea,
    input wire vga_bm0_wea,
    input wire vga_bt1_wea,
    input wire vga_bm1_wea,
    input wire vga_bmp_wea,
    input wire [23:0] cpu_addr,
    input wire [31:0] cpu_din,

    input wire cpu_reg_rd,
    output reg [31:0] cpu_dout,
    output reg cpu_ready,
    output reg cpu_hirq,
    output reg cpu_virq,

    // VGA signal Output
    output wire vga_hs,
    output wire vga_vs,
    output wire vga_blank,
    output reg [7:0] vga_r,
    output reg [7:0] vga_g,
    output reg [7:0] vga_b
    );

  // Video Registers

    // $000000 - Video Mode Bits - Default to BG0 Enabled Size:80x30 Scale:1x2 Pri:Highest, BG1 Disabled Size:64x64 Scale:2x2 Pri:Lowest
    reg [31:0] vid_mode = 32'b00000000110111000000100100000000;
    //      0 - Sprite Layer Enable
    //   7: 6 - Priority [00] Highest [11] Lowest
    //
    //      8 - BG Layer 0 Enable - 128x64
    //  10: 9 - Sizes: [00] 80x30, [01] 128x32, [10] 64x64, [11] 32x128
    //  13:11 - Scale: [000] 1x1, [001] 1x2, [010] 2x1, [011] 2x2, [100] 4x2, [101] 2x4, [110] 4x4, [111] 8x8
    //  15:14 - Priority [00] Highest [11] Lowest
    //
    //     16 - BG Layer 1 Enable - 128x64
    //  18:17 - Sizes: [00] 80x30, [01] 128x32, [10] 64x64, [11] 32x128
    //  21:19 - Scale: [000] 1x1, [001] 1x2, [010] 2x1, [011] 2x2, [100] 4x2, [101] 2x4, [110] 4x4, [111] 8x8
    //  23:22 - Priority [00] Highest [11] Lowest
    //
    //     24 - Bitmap Layer Enable - 256x128
    //  26:25 - Sizes: [00] 160x120, [01] 128x64, [10] 128x128, [11] 64x128
    //  29:27 - Scale: [000] 1x1, [001] 1x2, [010] 2x1, [011] 2x2, [100] 4x2, [101] 2x4, [110] 4x4, [111] 8x8
    //  31:30 - Priority [00] Highest [11] Lowest
    
    // $000020 - BG0 Scroll X (in Screen Pixels)
    reg [10:0] bg0_scroll_x = 0;
    // $000024 - BG0 Scroll Y (in Screen Pixels)
    reg [10:0] bg0_scroll_y = 0;
    // $000028 - BG0 Window X
    reg [31:0] bg0_window_x = 32'h02800000;
    wire [10:0] bg0_x1 = bg0_window_x[10:0];
    wire [10:0] bg0_x2 = bg0_window_x[26:16];
    // $00002C - BG0 Window Y
    reg [31:0] bg0_window_y = 32'h01B80028;
    wire [10:0] bg0_y1 = bg0_window_y[10:0];
    wire [10:0] bg0_y2 = bg0_window_y[26:16];
    // $000030 - BG0 Border Color
    reg [7:0] bg0_border = 8'h04;

    // $000040 - BG1 Scroll X (in Screen Pixels)
    reg [10:0] bg1_scroll_x = 0;
    // $000044 - BG1 Scroll Y (in Screen Pixels)
    reg [10:0] bg1_scroll_y = 0;
    // $000048 - BG1 Window X
    reg [31:0] bg1_window_x = 32'h02800000;
    wire [10:0] bg1_x1 = bg1_window_x[10:0];
    wire [10:0] bg1_x2 = bg1_window_x[26:16];
    // $00004C - BG1 Window Y
    reg [31:0] bg1_window_y = 32'h01E00000;
    wire [10:0] bg1_y1 = bg1_window_y[10:0];
    wire [10:0] bg1_y2 = bg1_window_y[26:16];
    // $000050 - BG1 Border Color
    reg [7:0] bg1_border = 8'h00;

    // $000060 - Bitmap Scroll X (in Screen Pixels)
    reg [10:0] bmp_scroll_x = 0;
    // $000064 - Bitmap Scroll Y (in Screen Pixels)
    reg [10:0] bmp_scroll_y = 0;
    // $000068 - Bitmap Window X
    reg [31:0] bmp_window_x = 32'h02800000;
    wire [10:0] bmp_x1 = bmp_window_x[10:0];
    wire [10:0] bmp_x2 = bmp_window_x[26:16];
    // $00006C - Bitmap Window Y
    reg [31:0] bmp_window_y = 32'h01E00000;
    wire [10:0] bmp_y1 = bmp_window_y[10:0];
    wire [10:0] bmp_y2 = bmp_window_y[26:16];
    // $000070 - Bitmap Border Color
    reg [7:0] bmp_border = 8'h00;

    //Horizontal
    // Sync is adjusted to compensate lower clock frequency
    reg [10:0] h_front   = 11'd40;  // 16;  // 18;  //Front porch
    reg [10:0] h_sync    = 11'd128; // 96;  // 96;  //Sync
    reg [10:0] h_back    = 11'd88;  // 48;  // 38;  //Back porch
    reg [10:0] h_active  = 11'd800; // 640; // 640; //Active pixels
    reg [10:0] h_irq     = 11'h2047; // Trigger H-Sync IRQ on this line at h_active

    //Vertical
    reg [10:0] v_front   = 11'd1;   // 10;  // 10;  //Front porch
    reg [10:0] v_sync    = 11'd4;   // 2;   // 2;   //Sync
    reg [10:0] v_back    = 11'd23;  // 33;  // 33;  //Back porch
    reg [10:0] v_active  = 11'd600; // 480; // 480; //Active lines // Trigger V-Sync IRQ on this line

    //X,Y positions generated by the timing generator
    wire [10:0] vga_x;
    wire [10:0] vga_y;

    always@(posedge cpu_clk) begin
        cpu_ready <= 1'b0;
        if (vga_reg_wea)
        begin
            case (cpu_addr[7:2])
                6'h00: vid_mode <= cpu_din[31:0];
                6'h01: begin
                    v_front <= cpu_din[26:16];
                    h_front <= cpu_din[10:0];
                end
                6'h02: begin
                    v_sync <= cpu_din[26:16];
                    h_sync <= cpu_din[10:0];
                end
                6'h03: begin
                    v_back <= cpu_din[26:16];
                    h_back <= cpu_din[10:0];
                end
                6'h04: begin
                    v_active <= cpu_din[26:16];
                    h_active <= cpu_din[10:0];
                end
                6'h05: begin
                    h_irq <= cpu_din[10:0];
                end
                6'h08: bg0_scroll_x <= cpu_din[10:0];
                6'h09: bg0_scroll_y <= cpu_din[10:0];
                6'h0A: bg0_window_x <= cpu_din[31:0];
                6'h0B: bg0_window_y <= cpu_din[31:0];
                6'h0C: bg0_border <= cpu_din[7:0];
                6'h10: bg1_scroll_x <= cpu_din[10:0];
                6'h11: bg1_scroll_y <= cpu_din[10:0];
                6'h12: bg1_window_x <= cpu_din[31:0];
                6'h13: bg1_window_y <= cpu_din[31:0];
                6'h14: bg1_border <= cpu_din[7:0];
                6'h18: bmp_scroll_x <= cpu_din[10:0];
                6'h19: bmp_scroll_y <= cpu_din[10:0];
                6'h1A: bmp_window_x <= cpu_din[31:0];
                6'h1B: bmp_window_y <= cpu_din[31:0];
                6'h1C: bmp_border <= cpu_din[7:0];
            endcase
            cpu_ready <= 1'b1;
        end
        if (cpu_reg_rd)
        begin
            case (cpu_addr[7:2])
               6'h00: cpu_dout <= vid_mode;
               6'h01: cpu_dout <= { 5'd0, v_front, 5'd0, h_front };
               6'h02: cpu_dout <= { 5'd0, v_sync, 5'd0, h_sync };
               6'h03: cpu_dout <= { 5'd0, v_back, 5'd0, h_back };
               6'h04: cpu_dout <= { 5'd0, v_active, 5'd0, h_active };
               6'h05: cpu_dout <= { 21'd0, vga_y };
               6'h08: cpu_dout <= { 21'd0, bg0_scroll_x };
               6'h09: cpu_dout <= { 21'd0, bg0_scroll_y };
               6'h0A: cpu_dout <= bg0_window_x;
               6'h0B: cpu_dout <= bg0_window_y;
               6'h0C: cpu_dout <= { 24'd0, bg0_border };
               6'h10: cpu_dout <= { 21'd0, bg1_scroll_x };
               6'h11: cpu_dout <= { 21'd0, bg1_scroll_y };
               6'h12: cpu_dout <= bg1_window_x;
               6'h13: cpu_dout <= bg1_window_y;
               6'h14: cpu_dout <= { 24'd0, bg1_border };
               6'h18: cpu_dout <= { 21'd0, bmp_scroll_x };
               6'h19: cpu_dout <= { 21'd0, bmp_scroll_y };
               6'h1A: cpu_dout <= bmp_window_x;
               6'h1B: cpu_dout <= bmp_window_y;
               6'h1C: cpu_dout <= { 24'd0, bmp_border };
            endcase        
            cpu_ready <= 1'b1;
        end
    end

    // Sprite Layer
    // Sprite Object Attribute Memory
    reg [31:0] spr_oam0_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam0_attr1 = 32'h00000000;
    reg [31:0] spr_oam1_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam1_attr1 = 32'h00000000;
    reg [31:0] spr_oam2_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam2_attr1 = 32'h00000000;
    reg [31:0] spr_oam3_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam3_attr1 = 32'h00000000;
    reg [31:0] spr_oam4_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam4_attr1 = 32'h00000000;
    reg [31:0] spr_oam5_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam5_attr1 = 32'h00000000;
    reg [31:0] spr_oam6_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam6_attr1 = 32'h00000000;
    reg [31:0] spr_oam7_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam7_attr1 = 32'h00000000;
    reg [31:0] spr_oam8_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam8_attr1 = 32'h00000000;
    reg [31:0] spr_oam9_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam9_attr1 = 32'h00000000;
    reg [31:0] spr_oam10_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam10_attr1 = 32'h00000000;
    reg [31:0] spr_oam11_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam11_attr1 = 32'h00000000;
    reg [31:0] spr_oam12_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam12_attr1 = 32'h00000000;
    reg [31:0] spr_oam13_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam13_attr1 = 32'h00000000;
    reg [31:0] spr_oam14_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam14_attr1 = 32'h00000000;
    reg [31:0] spr_oam15_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam15_attr1 = 32'h00000000;
    reg [31:0] spr_oam16_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam16_attr1 = 32'h00000000;
    reg [31:0] spr_oam17_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam17_attr1 = 32'h00000000;
    reg [31:0] spr_oam18_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam18_attr1 = 32'h00000000;
    reg [31:0] spr_oam19_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam19_attr1 = 32'h00000000;
    reg [31:0] spr_oam20_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam20_attr1 = 32'h00000000;
    reg [31:0] spr_oam21_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam21_attr1 = 32'h00000000;
    reg [31:0] spr_oam22_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam22_attr1 = 32'h00000000;
    reg [31:0] spr_oam23_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam23_attr1 = 32'h00000000;
    reg [31:0] spr_oam24_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam24_attr1 = 32'h00000000;
    reg [31:0] spr_oam25_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam25_attr1 = 32'h00000000;
    reg [31:0] spr_oam26_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam26_attr1 = 32'h00000000;
    reg [31:0] spr_oam27_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam27_attr1 = 32'h00000000;
    reg [31:0] spr_oam28_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam28_attr1 = 32'h00000000;
    reg [31:0] spr_oam29_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam29_attr1 = 32'h00000000;
    reg [31:0] spr_oam30_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam30_attr1 = 32'h00000000;
    reg [31:0] spr_oam31_attr0 = 32'hFFFFFFFF;
    reg [31:0] spr_oam31_attr1 = 32'h00000000;

    always@(posedge cpu_clk) begin
        if (vga_oam_wea)
        begin
            case (cpu_addr[7:2])
                6'h00: spr_oam0_attr0[31:0] <= cpu_din[31:0];
                6'h01: spr_oam0_attr1[31:0] <= cpu_din[31:0];
                6'h02: spr_oam1_attr0[31:0] <= cpu_din[31:0];
                6'h03: spr_oam1_attr1[31:0] <= cpu_din[31:0];
                6'h04: spr_oam2_attr0[31:0] <= cpu_din[31:0];
                6'h05: spr_oam2_attr1[31:0] <= cpu_din[31:0];
                6'h06: spr_oam3_attr0[31:0] <= cpu_din[31:0];
                6'h07: spr_oam3_attr1[31:0] <= cpu_din[31:0];
                6'h08: spr_oam4_attr0[31:0] <= cpu_din[31:0];
                6'h09: spr_oam4_attr1[31:0] <= cpu_din[31:0];
                6'h0A: spr_oam5_attr0[31:0] <= cpu_din[31:0];
                6'h0B: spr_oam5_attr1[31:0] <= cpu_din[31:0];
                6'h0C: spr_oam6_attr0[31:0] <= cpu_din[31:0];
                6'h0D: spr_oam6_attr1[31:0] <= cpu_din[31:0];
                6'h0E: spr_oam7_attr0[31:0] <= cpu_din[31:0];
                6'h0F: spr_oam7_attr1[31:0] <= cpu_din[31:0];
                6'h10: spr_oam8_attr0[31:0] <= cpu_din[31:0];
                6'h11: spr_oam8_attr1[31:0] <= cpu_din[31:0];
                6'h12: spr_oam9_attr0[31:0] <= cpu_din[31:0];
                6'h13: spr_oam9_attr1[31:0] <= cpu_din[31:0];
                6'h14: spr_oam10_attr0[31:0] <= cpu_din[31:0];
                6'h15: spr_oam10_attr1[31:0] <= cpu_din[31:0];
                6'h16: spr_oam11_attr0[31:0] <= cpu_din[31:0];
                6'h17: spr_oam11_attr1[31:0] <= cpu_din[31:0];
                6'h18: spr_oam12_attr0[31:0] <= cpu_din[31:0];
                6'h19: spr_oam12_attr1[31:0] <= cpu_din[31:0];
                6'h1A: spr_oam13_attr0[31:0] <= cpu_din[31:0];
                6'h1B: spr_oam13_attr1[31:0] <= cpu_din[31:0];
                6'h1C: spr_oam14_attr0[31:0] <= cpu_din[31:0];
                6'h1D: spr_oam14_attr1[31:0] <= cpu_din[31:0];
                6'h1E: spr_oam15_attr0[31:0] <= cpu_din[31:0];
                6'h1F: spr_oam15_attr1[31:0] <= cpu_din[31:0];
                6'h20: spr_oam16_attr0[31:0] <= cpu_din[31:0];
                6'h21: spr_oam16_attr1[31:0] <= cpu_din[31:0];
                6'h22: spr_oam17_attr0[31:0] <= cpu_din[31:0];
                6'h23: spr_oam17_attr1[31:0] <= cpu_din[31:0];
                6'h24: spr_oam18_attr0[31:0] <= cpu_din[31:0];
                6'h25: spr_oam18_attr1[31:0] <= cpu_din[31:0];
                6'h26: spr_oam19_attr0[31:0] <= cpu_din[31:0];
                6'h27: spr_oam19_attr1[31:0] <= cpu_din[31:0];
                6'h28: spr_oam20_attr0[31:0] <= cpu_din[31:0];
                6'h29: spr_oam20_attr1[31:0] <= cpu_din[31:0];
                6'h2A: spr_oam21_attr0[31:0] <= cpu_din[31:0];
                6'h2B: spr_oam21_attr1[31:0] <= cpu_din[31:0];
                6'h2C: spr_oam22_attr0[31:0] <= cpu_din[31:0];
                6'h2D: spr_oam22_attr1[31:0] <= cpu_din[31:0];
                6'h2E: spr_oam23_attr0[31:0] <= cpu_din[31:0];
                6'h2F: spr_oam23_attr1[31:0] <= cpu_din[31:0];
                6'h30: spr_oam24_attr0[31:0] <= cpu_din[31:0];
                6'h31: spr_oam24_attr1[31:0] <= cpu_din[31:0];
                6'h32: spr_oam25_attr0[31:0] <= cpu_din[31:0];
                6'h33: spr_oam25_attr1[31:0] <= cpu_din[31:0];
                6'h34: spr_oam26_attr0[31:0] <= cpu_din[31:0];
                6'h35: spr_oam26_attr1[31:0] <= cpu_din[31:0];
                6'h36: spr_oam27_attr0[31:0] <= cpu_din[31:0];
                6'h37: spr_oam27_attr1[31:0] <= cpu_din[31:0];
                6'h38: spr_oam28_attr0[31:0] <= cpu_din[31:0];
                6'h39: spr_oam28_attr1[31:0] <= cpu_din[31:0];
                6'h3A: spr_oam29_attr0[31:0] <= cpu_din[31:0];
                6'h3B: spr_oam29_attr1[31:0] <= cpu_din[31:0];
                6'h3C: spr_oam30_attr0[31:0] <= cpu_din[31:0];
                6'h3D: spr_oam30_attr1[31:0] <= cpu_din[31:0];
                6'h3E: spr_oam31_attr0[31:0] <= cpu_din[31:0];
                6'h3F: spr_oam31_attr1[31:0] <= cpu_din[31:0];
            endcase
        end
    end

    wire sprite0_visible;
    wire [14:0] sprite0_tile_addr;
    wire [3:0] sprite0_pal;
    sprite sprite0(
        .vga_clk(!vga_clk),
        .attr0(spr_oam0_attr0[31:0]),
        .attr1(spr_oam0_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite0_tile_addr[14:0]),
        .spr_pal(sprite0_pal[3:0]),
        .visible(sprite0_visible)
    );
    wire sprite1_visible;
    wire [14:0] sprite1_tile_addr;
    wire [3:0] sprite1_pal;
    sprite sprite1(
        .vga_clk(vga_clk),
        .attr0(spr_oam1_attr0[31:0]),
        .attr1(spr_oam1_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite1_tile_addr[14:0]),
        .spr_pal(sprite1_pal[3:0]),
        .visible(sprite1_visible)
    );
    wire sprite2_visible;
    wire [14:0] sprite2_tile_addr;
    wire [3:0] sprite2_pal;
    sprite sprite2(
        .vga_clk(vga_clk),
        .attr0(spr_oam2_attr0[31:0]),
        .attr1(spr_oam2_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite2_tile_addr[14:0]),
        .spr_pal(sprite2_pal[3:0]),
        .visible(sprite2_visible)
    );
    wire sprite3_visible;
    wire [14:0] sprite3_tile_addr;
    wire [3:0] sprite3_pal;
    sprite sprite3(
        .vga_clk(vga_clk),
        .attr0(spr_oam3_attr0[31:0]),
        .attr1(spr_oam3_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite3_tile_addr[14:0]),
        .spr_pal(sprite3_pal[3:0]),
        .visible(sprite3_visible)
    );
    wire sprite4_visible;
    wire [14:0] sprite4_tile_addr;
    wire [3:0] sprite4_pal;
    sprite sprite4(
        .vga_clk(!vga_clk),
        .attr0(spr_oam4_attr0[31:0]),
        .attr1(spr_oam4_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite4_tile_addr[14:0]),
        .spr_pal(sprite4_pal[3:0]),
        .visible(sprite4_visible)
    );
    wire sprite5_visible;
    wire [14:0] sprite5_tile_addr;
    wire [3:0] sprite5_pal;
    sprite sprite5(
        .vga_clk(vga_clk),
        .attr0(spr_oam5_attr0[31:0]),
        .attr1(spr_oam5_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite5_tile_addr[14:0]),
        .spr_pal(sprite5_pal[3:0]),
        .visible(sprite5_visible)
    );
    wire sprite6_visible;
    wire [14:0] sprite6_tile_addr;
    wire [3:0] sprite6_pal;
    sprite sprite6(
        .vga_clk(vga_clk),
        .attr0(spr_oam6_attr0[31:0]),
        .attr1(spr_oam6_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite6_tile_addr[14:0]),
        .spr_pal(sprite6_pal[3:0]),
        .visible(sprite6_visible)
    );
    wire sprite7_visible;
    wire [14:0] sprite7_tile_addr;
    wire [3:0] sprite7_pal;
    sprite sprite7(
        .vga_clk(vga_clk),
        .attr0(spr_oam7_attr0[31:0]),
        .attr1(spr_oam7_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite7_tile_addr[14:0]),
        .spr_pal(sprite7_pal[3:0]),
        .visible(sprite7_visible)
    );
    wire sprite8_visible;
    wire [14:0] sprite8_tile_addr;
    wire [3:0] sprite8_pal;
    sprite sprite8(
        .vga_clk(!vga_clk),
        .attr0(spr_oam8_attr0[31:0]),
        .attr1(spr_oam8_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite8_tile_addr[14:0]),
        .spr_pal(sprite8_pal[3:0]),
        .visible(sprite8_visible)
    );
    wire sprite9_visible;
    wire [14:0] sprite9_tile_addr;
    wire [3:0] sprite9_pal;
    sprite sprite9(
        .vga_clk(vga_clk),
        .attr0(spr_oam9_attr0[31:0]),
        .attr1(spr_oam9_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite9_tile_addr[14:0]),
        .spr_pal(sprite9_pal[3:0]),
        .visible(sprite9_visible)
    );
    wire sprite10_visible;
    wire [14:0] sprite10_tile_addr;
    wire [3:0] sprite10_pal;
    sprite sprite10(
        .vga_clk(vga_clk),
        .attr0(spr_oam10_attr0[31:0]),
        .attr1(spr_oam10_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite10_tile_addr[14:0]),
        .spr_pal(sprite10_pal[3:0]),
        .visible(sprite10_visible)
    );
    wire sprite11_visible;
    wire [14:0] sprite11_tile_addr;
    wire [3:0] sprite11_pal;
    sprite sprite11(
        .vga_clk(vga_clk),
        .attr0(spr_oam11_attr0[31:0]),
        .attr1(spr_oam11_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite11_tile_addr[14:0]),
        .spr_pal(sprite11_pal[3:0]),
        .visible(sprite11_visible)
    );
    wire sprite12_visible;
    wire [14:0] sprite12_tile_addr;
    wire [3:0] sprite12_pal;
    sprite sprite12(
        .vga_clk(!vga_clk),
        .attr0(spr_oam12_attr0[31:0]),
        .attr1(spr_oam12_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite12_tile_addr[14:0]),
        .spr_pal(sprite12_pal[3:0]),
        .visible(sprite12_visible)
    );
    wire sprite13_visible;
    wire [14:0] sprite13_tile_addr;
    wire [3:0] sprite13_pal;
    sprite sprite13(
        .vga_clk(vga_clk),
        .attr0(spr_oam13_attr0[31:0]),
        .attr1(spr_oam13_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite13_tile_addr[14:0]),
        .spr_pal(sprite13_pal[3:0]),
        .visible(sprite13_visible)
    );
    wire sprite14_visible;
    wire [14:0] sprite14_tile_addr;
    wire [3:0] sprite14_pal;
    sprite sprite14(
        .vga_clk(vga_clk),
        .attr0(spr_oam14_attr0[31:0]),
        .attr1(spr_oam14_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite14_tile_addr[14:0]),
        .spr_pal(sprite14_pal[3:0]),
        .visible(sprite14_visible)
    );
    wire sprite15_visible;
    wire [14:0] sprite15_tile_addr;
    wire [3:0] sprite15_pal;
    sprite sprite15(
        .vga_clk(vga_clk),
        .attr0(spr_oam15_attr0[31:0]),
        .attr1(spr_oam15_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite15_tile_addr[14:0]),
        .spr_pal(sprite15_pal[3:0]),
        .visible(sprite15_visible)
    );
    wire sprite16_visible;
    wire [14:0] sprite16_tile_addr;
    wire [3:0] sprite16_pal;
    sprite sprite16(
        .vga_clk(vga_clk),
        .attr0(spr_oam16_attr0[31:0]),
        .attr1(spr_oam16_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite16_tile_addr[14:0]),
        .spr_pal(sprite16_pal[3:0]),
        .visible(sprite16_visible)
    );
    wire sprite17_visible;
    wire [14:0] sprite17_tile_addr;
    wire [3:0] sprite17_pal;
    sprite sprite17(
        .vga_clk(vga_clk),
        .attr0(spr_oam17_attr0[31:0]),
        .attr1(spr_oam17_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite17_tile_addr[14:0]),
        .spr_pal(sprite17_pal[3:0]),
        .visible(sprite17_visible)
    );
    wire sprite18_visible;
    wire [14:0] sprite18_tile_addr;
    wire [3:0] sprite18_pal;
    sprite sprite18(
        .vga_clk(!vga_clk),
        .attr0(spr_oam18_attr0[31:0]),
        .attr1(spr_oam18_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite18_tile_addr[14:0]),
        .spr_pal(sprite18_pal[3:0]),
        .visible(sprite18_visible)
    );
    wire sprite19_visible;
    wire [14:0] sprite19_tile_addr;
    wire [3:0] sprite19_pal;
    sprite sprite19(
        .vga_clk(vga_clk),
        .attr0(spr_oam19_attr0[31:0]),
        .attr1(spr_oam19_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite19_tile_addr[14:0]),
        .spr_pal(sprite19_pal[3:0]),
        .visible(sprite19_visible)
    );
    wire sprite20_visible;
    wire [14:0] sprite20_tile_addr;
    wire [3:0] sprite20_pal;
    sprite sprite20(
        .vga_clk(!vga_clk),
        .attr0(spr_oam20_attr0[31:0]),
        .attr1(spr_oam20_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite20_tile_addr[14:0]),
        .spr_pal(sprite20_pal[3:0]),
        .visible(sprite20_visible)
    );
    wire sprite21_visible;
    wire [14:0] sprite21_tile_addr;
    wire [3:0] sprite21_pal;
    sprite sprite21(
        .vga_clk(vga_clk),
        .attr0(spr_oam21_attr0[31:0]),
        .attr1(spr_oam21_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite21_tile_addr[14:0]),
        .spr_pal(sprite21_pal[3:0]),
        .visible(sprite21_visible)
    );
    wire sprite22_visible;
    wire [14:0] sprite22_tile_addr;
    wire [3:0] sprite22_pal;
    sprite sprite22(
        .vga_clk(vga_clk),
        .attr0(spr_oam22_attr0[31:0]),
        .attr1(spr_oam22_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite22_tile_addr[14:0]),
        .spr_pal(sprite22_pal[3:0]),
        .visible(sprite22_visible)
    );
    wire sprite23_visible;
    wire [14:0] sprite23_tile_addr;
    wire [3:0] sprite23_pal;
    sprite sprite23(
        .vga_clk(vga_clk),
        .attr0(spr_oam23_attr0[31:0]),
        .attr1(spr_oam23_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite23_tile_addr[14:0]),
        .spr_pal(sprite23_pal[3:0]),
        .visible(sprite23_visible)
    );
    wire sprite24_visible;
    wire [14:0] sprite24_tile_addr;
    wire [3:0] sprite24_pal;
    sprite sprite24(
        .vga_clk(!vga_clk),
        .attr0(spr_oam24_attr0[31:0]),
        .attr1(spr_oam24_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite24_tile_addr[14:0]),
        .spr_pal(sprite24_pal[3:0]),
        .visible(sprite24_visible)
    );
    wire sprite25_visible;
    wire [14:0] sprite25_tile_addr;
    wire [3:0] sprite25_pal;
    sprite sprite25(
        .vga_clk(vga_clk),
        .attr0(spr_oam25_attr0[31:0]),
        .attr1(spr_oam25_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite25_tile_addr[14:0]),
        .spr_pal(sprite25_pal[3:0]),
        .visible(sprite25_visible)
    );
    wire sprite26_visible;
    wire [14:0] sprite26_tile_addr;
    wire [3:0] sprite26_pal;
    sprite sprite26(
        .vga_clk(vga_clk),
        .attr0(spr_oam26_attr0[31:0]),
        .attr1(spr_oam26_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite26_tile_addr[14:0]),
        .spr_pal(sprite26_pal[3:0]),
        .visible(sprite26_visible)
    );
    wire sprite27_visible;
    wire [14:0] sprite27_tile_addr;
    wire [3:0] sprite27_pal;
    sprite sprite27(
        .vga_clk(vga_clk),
        .attr0(spr_oam27_attr0[31:0]),
        .attr1(spr_oam27_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite27_tile_addr[14:0]),
        .spr_pal(sprite27_pal[3:0]),
        .visible(sprite27_visible)
    );
    wire sprite28_visible;
    wire [14:0] sprite28_tile_addr;
    wire [3:0] sprite28_pal;
    sprite sprite28(
        .vga_clk(!vga_clk),
        .attr0(spr_oam28_attr0[31:0]),
        .attr1(spr_oam28_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite28_tile_addr[14:0]),
        .spr_pal(sprite28_pal[3:0]),
        .visible(sprite28_visible)
    );
    wire sprite29_visible;
    wire [14:0] sprite29_tile_addr;
    wire [3:0] sprite29_pal;
    sprite sprite29(
        .vga_clk(vga_clk),
        .attr0(spr_oam29_attr0[31:0]),
        .attr1(spr_oam29_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite29_tile_addr[14:0]),
        .spr_pal(sprite29_pal[3:0]),
        .visible(sprite29_visible)
    );
    wire sprite30_visible;
    wire [14:0] sprite30_tile_addr;
    wire [3:0] sprite30_pal;
    sprite sprite30(
        .vga_clk(vga_clk),
        .attr0(spr_oam30_attr0[31:0]),
        .attr1(spr_oam30_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite30_tile_addr[14:0]),
        .spr_pal(sprite30_pal[3:0]),
        .visible(sprite30_visible)
    );
    wire sprite31_visible;
    wire [14:0] sprite31_tile_addr;
    wire [3:0] sprite31_pal;
    sprite sprite31(
        .vga_clk(vga_clk),
        .attr0(spr_oam31_attr0[31:0]),
        .attr1(spr_oam31_attr1[31:0]),
        .vga_x(vga_x[10:0]),
        .vga_y(vga_y[10:0]),
        .tile_addr(sprite31_tile_addr[14:0]),
        .spr_pal(sprite31_pal[3:0]),
        .visible(sprite31_visible)
    );
    
    // Sprite Map is 4-Bits per Pixel
    wire spr_enable = vid_mode[0];
    wire [1:0] spr_priority = vid_mode[7:6];
    wire spr_active = spr_enable & (
        sprite0_visible | sprite1_visible | sprite2_visible | sprite3_visible | sprite4_visible | sprite5_visible | sprite6_visible | sprite7_visible |
        sprite8_visible | sprite9_visible | sprite10_visible | sprite11_visible | sprite12_visible | sprite13_visible | sprite14_visible | sprite15_visible |
        sprite16_visible | sprite17_visible | sprite18_visible | sprite19_visible | sprite20_visible | sprite21_visible | sprite22_visible | sprite23_visible |
        sprite24_visible | sprite25_visible | sprite26_visible | sprite27_visible | sprite28_visible | sprite29_visible | sprite30_visible | sprite31_visible
        );
    wire [3:0] spr_map_dout;
    wire [14:0] spr_map_addr = 
        ((sprite0_visible) ? sprite0_tile_addr[14:0] : 
        ((sprite1_visible) ? sprite1_tile_addr[14:0] : 
        ((sprite2_visible) ? sprite2_tile_addr[14:0] : 
        ((sprite3_visible) ? sprite3_tile_addr[14:0] : 
        ((sprite4_visible) ? sprite4_tile_addr[14:0] : 
        ((sprite5_visible) ? sprite5_tile_addr[14:0] : 
        ((sprite6_visible) ? sprite6_tile_addr[14:0] : 
        ((sprite7_visible) ? sprite7_tile_addr[14:0] : 
        ((sprite8_visible) ? sprite8_tile_addr[14:0] : 
        ((sprite9_visible) ? sprite9_tile_addr[14:0] : 
        ((sprite10_visible) ? sprite10_tile_addr[14:0] : 
        ((sprite11_visible) ? sprite11_tile_addr[14:0] : 
        ((sprite12_visible) ? sprite12_tile_addr[14:0] : 
        ((sprite13_visible) ? sprite13_tile_addr[14:0] : 
        ((sprite14_visible) ? sprite14_tile_addr[14:0] : 
        ((sprite15_visible) ? sprite15_tile_addr[14:0] : 
        ((sprite16_visible) ? sprite16_tile_addr[14:0] : 
        ((sprite17_visible) ? sprite17_tile_addr[14:0] : 
        ((sprite18_visible) ? sprite18_tile_addr[14:0] : 
        ((sprite19_visible) ? sprite19_tile_addr[14:0] : 
        ((sprite20_visible) ? sprite20_tile_addr[14:0] : 
        ((sprite21_visible) ? sprite21_tile_addr[14:0] : 
        ((sprite22_visible) ? sprite22_tile_addr[14:0] : 
        ((sprite23_visible) ? sprite23_tile_addr[14:0] : 
        ((sprite24_visible) ? sprite24_tile_addr[14:0] : 
        ((sprite25_visible) ? sprite25_tile_addr[14:0] : 
        ((sprite26_visible) ? sprite26_tile_addr[14:0] : 
        ((sprite27_visible) ? sprite27_tile_addr[14:0] : 
        ((sprite28_visible) ? sprite28_tile_addr[14:0] : 
        ((sprite29_visible) ? sprite29_tile_addr[14:0] : 
        ((sprite30_visible) ? sprite30_tile_addr[14:0] : 
        ((sprite31_visible) ? sprite31_tile_addr[14:0] : 
        0))))))))))))))))))))))))))))))));
    wire [3:0] spr_palidx = 
        ((sprite0_visible) ? sprite0_pal[3:0] : 
        ((sprite1_visible) ? sprite1_pal[3:0] : 
        ((sprite2_visible) ? sprite2_pal[3:0] : 
        ((sprite3_visible) ? sprite3_pal[3:0] : 
        ((sprite4_visible) ? sprite4_pal[3:0] : 
        ((sprite5_visible) ? sprite5_pal[3:0] : 
        ((sprite6_visible) ? sprite6_pal[3:0] : 
        ((sprite7_visible) ? sprite7_pal[3:0] : 
        ((sprite8_visible) ? sprite8_pal[3:0] : 
        ((sprite9_visible) ? sprite9_pal[3:0] : 
        ((sprite10_visible) ? sprite10_pal[3:0] : 
        ((sprite11_visible) ? sprite11_pal[3:0] : 
        ((sprite12_visible) ? sprite12_pal[3:0] : 
        ((sprite13_visible) ? sprite13_pal[3:0] : 
        ((sprite14_visible) ? sprite14_pal[3:0] : 
        ((sprite15_visible) ? sprite15_pal[3:0] : 
        ((sprite16_visible) ? sprite16_pal[3:0] : 
        ((sprite17_visible) ? sprite17_pal[3:0] : 
        ((sprite18_visible) ? sprite18_pal[3:0] : 
        ((sprite19_visible) ? sprite19_pal[3:0] : 
        ((sprite20_visible) ? sprite20_pal[3:0] : 
        ((sprite21_visible) ? sprite21_pal[3:0] : 
        ((sprite22_visible) ? sprite22_pal[3:0] : 
        ((sprite23_visible) ? sprite23_pal[3:0] : 
        ((sprite24_visible) ? sprite24_pal[3:0] : 
        ((sprite25_visible) ? sprite25_pal[3:0] : 
        ((sprite26_visible) ? sprite26_pal[3:0] : 
        ((sprite27_visible) ? sprite27_pal[3:0] : 
        ((sprite28_visible) ? sprite28_pal[3:0] : 
        ((sprite29_visible) ? sprite29_pal[3:0] : 
        ((sprite30_visible) ? sprite30_pal[3:0] : 
        ((sprite31_visible) ? sprite31_pal[3:0] : 
        0))))))))))))))))))))))))))))))));
    spr_map spr_map(
        .clka(!cpu_clk),
        .wea(vga_spr_wea),
        .addra(cpu_addr[16:2]),
        .dina(cpu_din[3:0]),
        .clkb(vga_clk),
        .addrb(spr_map_addr[14:0]),
        .doutb(spr_map_dout)
    );
    wire [7:0] spr_color = ((spr_active) && (spr_map_dout[3:0] != 4'd0)) ? ( (spr_palidx[3:0] << 4) | spr_map_dout[3:0] ) : 8'h00;


    // BG Layer 0 is 24-bit wide 180x30 (normally used for 80x25, 80x30, 40x25, 40x30 Text)
    //   6:0  - Tile Index
    //  15:8  - BG color
    //  23:16 - FG color
    // BG0 Map is 1-Bit per Pixel
    wire bg0_enable = vid_mode[8];
    wire [1:0] bg0_size = vid_mode[10:9];
    wire [2:0] bg0_scale = vid_mode[13:11];
    wire bg0_active = (bg0_enable) && (vga_x[10:0] >= bg0_x1[10:0]) && (vga_x[10:0] <= bg0_x2[10:0]) && (vga_y[10:0] >= bg0_y1[10:0]) && (vga_y[10:0] <= bg0_y2[10:0]);
    wire [1:0] bg0_priority = vid_mode[15:14];
    wire [10:0] bg0_xx = (vga_x[10:0] - bg0_scroll_x[10:0]);
    wire [9:0] bg0_x =
        ((bg0_scale[2:0] == 3'b111) ? (bg0_xx[10:3]) :
        ((bg0_scale[2:0] == 3'b110) ? (bg0_xx[10:2]) :
        ((bg0_scale[2:0] == 3'b101) ? (bg0_xx[10:1]) :
        ((bg0_scale[2:0] == 3'b100) ? (bg0_xx[10:1]) :
        ((bg0_scale[2:0] == 3'b010) ? (bg0_xx[10:1]) :
        ((bg0_scale[2:0] == 3'b011) ? (bg0_xx[10:1]) :
        (bg0_xx[10:0])))))));
    wire [10:0] bg0_yy = (vga_y[10:0] - bg0_scroll_y[10:0]);
    wire [9:0] bg0_y =
        ((bg0_scale[2:0] == 3'b111) ? (bg0_yy[10:3]) :
        ((bg0_scale[2:0] == 3'b101) ? (bg0_yy[10:2]) :
        ((bg0_scale[2:0] == 3'b110) ? (bg0_yy[10:1]) :
        ((bg0_scale[2:0] == 3'b100) ? (bg0_yy[10:1]) :
        ((bg0_scale[2:0] == 3'b001) ? (bg0_yy[10:1]) :
        ((bg0_scale[2:0] == 3'b011) ? (bg0_yy[10:1]) :
        (bg0_yy[10:0])))))));
    wire [6:0] bg0_tile_x = bg0_x[9:3];
    wire [6:0] bg0_tile_y = bg0_y[9:3];
    wire [11:0] bg0_til_addr = 
        ((bg0_size == 2'b00) ? (bg0_tile_y[5:0] * 80 + bg0_tile_x[6:0]) :
        ((bg0_size == 2'b01) ? ((bg0_tile_y[4:0] << 7) | bg0_tile_x[6:0]) :
        ((bg0_size == 2'b10) ? ((bg0_tile_y[5:0] << 6) | bg0_tile_x[5:0]) :
        /*(bg0_size == 2'b11) ?*/ ((bg0_tile_y[6:0] << 5) | bg0_tile_x[4:0]))));
    wire [23:0] bg0_til_dout;
    bg0_til bg0_til(
        .clka(!cpu_clk),
        .wea(vga_bt0_wea),
        .addra(cpu_addr[13:2]),
        .dina(cpu_din[23:0]),
        .clkb(!vga_clk),
        .addrb(bg0_til_addr[11:0]),
        .doutb(bg0_til_dout)
    );
    wire [7:0] bg0_tile = bg0_til_dout[7:0];
    wire [7:0] bg0_fg_color = bg0_til_dout[23:16];
    wire [7:0] bg0_bg_color = bg0_til_dout[15:8];

    //{ascii_code[7:1], ~ascii_code[0], row, ~col}
    //{bg0_tile[7:1], ~bg0_tile[0], ~bg0_y[2:0], ~bg0_x[2:0]}; //
    wire [13:0] bg0_map_addr = (bg0_tile << 6) | (bg0_y[2:0] << 3) | bg0_x[2:0];
    wire bg0_map_dout;
    bg0_map bg0_map(
        .clka(!cpu_clk),
        .wea(vga_bm0_wea),
        .addra(cpu_addr[15:2]),
        .dina(cpu_din[0]),
        .clkb(vga_clk),
        .addrb(bg0_map_addr[13:0]),
        .doutb(bg0_map_dout)
    );
    wire [7:0] bg0_color = (bg0_active) ? ((bg0_map_dout) ? (bg0_fg_color[7:0]) : (bg0_bg_color[7:0])) : bg0_border[7:0];


    // BG Layer 1 is 16-bit wide 128x64
    //   9:0  - Tile Index
    //   10   - H-Flip
    //   11   - V-Flip
    //  15:12 - Palette Hi Nybble
    // BG1 Map is 4-Bits per Pixel, providing the Low Nybble
    wire bg1_enable = vid_mode[16];
    wire [1:0] bg1_size = vid_mode[18:17];
    wire [2:0] bg1_scale = vid_mode[21:19];
    wire bg1_active = (bg1_enable) && (vga_x[10:0] >= bg1_x1[10:0]) && (vga_x[10:0] <= bg1_x2[10:0]) && (vga_y[10:0] >= bg1_y1[10:0]) && (vga_y[10:0] <= bg1_y2[10:0]);
    wire [1:0] bg1_priority = vid_mode[23:22];
    wire [10:0] bg1_xx = (vga_x - bg1_scroll_x);
    wire [9:0] bg1_x =
        ((bg1_scale[2:0] == 3'b111) ? (bg1_xx >> 3) :
        ((bg1_scale[2:0] == 3'b110) ? (bg1_xx >> 2) :
        ((bg1_scale[2:0] == 3'b101) ? (bg1_xx >> 1) :
        ((bg1_scale[2:0] == 3'b100) ? (bg1_xx >> 1) :
        ((bg1_scale[2:0] == 3'b010) ? (bg1_xx >> 1) :
        ((bg1_scale[2:0] == 3'b011) ? (bg1_xx >> 1) :
        (bg1_xx)))))));
    wire [10:0] bg1_yy = (vga_y - bg1_scroll_y);
    wire [9:0] bg1_y =
        ((bg1_scale[2:0] == 3'b111) ? (bg1_yy >> 3) :
        ((bg1_scale[2:0] == 3'b101) ? (bg1_yy >> 2) :
        ((bg1_scale[2:0] == 3'b110) ? (bg1_yy >> 1) :
        ((bg1_scale[2:0] == 3'b100) ? (bg1_yy >> 1) :
        ((bg1_scale[2:0] == 3'b001) ? (bg1_yy >> 1) :
        ((bg1_scale[2:0] == 3'b011) ? (bg1_yy >> 1) :
        (bg1_yy)))))));
    wire [6:0] bg1_tile_x = bg1_x[9:3];
    wire [6:0] bg1_tile_y = bg1_y[8:3];
    wire [12:0] bg1_til_addr = 
        ((bg1_size == 2'b00) ? (bg1_tile_y[5:0] * 80 + bg1_tile_x[6:0]) :
        ((bg1_size == 2'b01) ? ((bg1_tile_y[4:0] << 7) | bg1_tile_x[6:0]) :
        ((bg1_size == 2'b10) ? ((bg1_tile_y[5:0] << 6) | bg1_tile_x[5:0]) :
        /*(bg0_size == 2'b11) ?*/ ((bg1_tile_y[6:0] << 5) | bg1_tile_x[4:0]))));
    wire [15:0] bg1_til_dout;
    bg1_til bg1_til(
        .clka(!cpu_clk),
        .wea(vga_bt1_wea),
        .addra(cpu_addr[14:2]),
        .dina(cpu_din[23:0]),
        .clkb(!vga_clk),
        .addrb(bg1_til_addr[12:0]),
        .doutb(bg1_til_dout)
    );
    wire [9:0] bg1_tile = bg1_til_dout[9:0];
    wire bg1_flipx = bg1_til_dout[10];
    wire bg1_flipy = bg1_til_dout[11];
    wire [3:0] bg1_palidx = bg1_til_dout[15:12];

    wire [3:0] bg1_map_dout;
    wire [15:0] bg1_map_addr = (bg1_tile << 6) | (((bg1_flipy) ? (7 - bg1_y[2:0]) : bg1_y[2:0]) << 3) | ((bg1_flipx) ? (7 - bg1_x[2:0]) : bg1_x[2:0]);
    bg1_map bg1_map(
        .clka(!cpu_clk),
        .wea(vga_bm1_wea),
        .addra(cpu_addr[15:2]),
        .dina(cpu_din[3:0]),
        .clkb(vga_clk),
        .addrb(bg1_map_addr[13:0]),
        .doutb(bg1_map_dout)
    );
    wire [7:0] bg1_color = (bg1_active) ? ((bg1_palidx[3:0] << 4) | bg1_map_dout[3:0]) : bg1_border[7:0];

    
    // Bitmap Layer
    wire bmp_enable = vid_mode[24];
    wire [2:0] bmp_scale = vid_mode[27:25];
    wire bmp_active = bmp_enable & (vga_x >= bmp_x1) & (vga_x <= bmp_x2) & (vga_y >= bmp_y1) & (vga_y <= bmp_y2);
    wire [1:0] bmp_priority = vid_mode[31:30];
    wire [10:0] bmp_xx = (vga_x - bmp_scroll_x);
    wire [9:0] bmp_x =
        ((bmp_scale[2:0] == 3'b111) ? (bmp_xx >> 3) :
        ((bmp_scale[2:0] == 3'b110) ? (bmp_xx >> 2) :
        ((bmp_scale[2:0] == 3'b101) ? (bmp_xx >> 1) :
        ((bmp_scale[2:0] == 3'b100) ? (bmp_xx >> 1) :
        ((bmp_scale[2:0] == 3'b010) ? (bmp_xx >> 1) :
        ((bmp_scale[2:0] == 3'b011) ? (bmp_xx >> 1) :
        (bg1_xx)))))));
    wire [10:0] bmp_yy = (vga_y - bmp_scroll_y);
    wire [9:0] bmp_y =
        ((bmp_scale[2:0] == 3'b111) ? (bmp_yy >> 3) :
        ((bmp_scale[2:0] == 3'b101) ? (bmp_yy >> 2) :
        ((bmp_scale[2:0] == 3'b110) ? (bmp_yy >> 1) :
        ((bmp_scale[2:0] == 3'b100) ? (bmp_yy >> 1) :
        ((bmp_scale[2:0] == 3'b001) ? (bmp_yy >> 1) :
        ((bmp_scale[2:0] == 3'b011) ? (bmp_yy >> 1) :
        (bmp_yy)))))));
    wire [7:0] bmpcop_dout;
    wire [14:0] bmp_addr = bmp_y * 256 + bmp_x;
    copper_ram bmpcop(
        .clka(cpu_clk),
        .wea(vga_cop_wea),
        .addra(cpu_addr[12:2]),
        .dina(cpu_din[7:0]),
        .clkb(vga_clk),
        .addrb(bmp_yy[10:0]),
        .doutb(bmpcop_dout)
    );
    wire [1:0] bmpram_dout;
    bitmap_ram bmpram(
        .clka(cpu_clk),
        .wea(vga_bmp_wea),
        .addra(cpu_addr[16:2]),
        .dina(cpu_din[7:0]),
        .clkb(!vga_clk),
        .addrb(bmp_addr),
        .doutb(bmpram_dout)
    );
    wire [7:0] bmp_color = bmpcop_dout[7:0] + bmpram_dout[1:0];
    
    
    // Palette Lookup
    wire [7:0] pixel_lut = 
    
           // Priority 0
           (((bmp_priority[1:0] == 2'd0) && (bmp_color[7:0] != 8'h00)) ? bmp_color[7:0] :
           (((bg1_priority[1:0] == 2'd0) && (bg1_color[7:0] != 8'h00)) ? bg1_color[7:0] :
           (((bg0_priority[1:0] == 2'd0) && (bg0_color[7:0] != 8'h00)) ? bg0_color[7:0] :
           (((spr_priority[1:0] == 2'd0) && (spr_color[7:0] != 8'h00)) ? spr_color[7:0] :

           // Priority 1
           (((bmp_priority[1:0] == 2'd1) && (bmp_color[7:0] != 8'h00)) ? bmp_color[7:0] :
           (((bg1_priority[1:0] == 2'd1) && (bg1_color[7:0] != 8'h00)) ? bg1_color[7:0] :
           (((bg0_priority[1:0] == 2'd1) && (bg0_color[7:0] != 8'h00)) ? bg0_color[7:0] :
           (((spr_priority[1:0] == 2'd1) && (spr_color[7:0] != 8'h00)) ? spr_color[7:0] :

           // Priority 2
           (((bmp_priority[1:0] == 2'd2) && (bmp_color[7:0] != 8'h00)) ? bmp_color[7:0] :
           (((bg1_priority[1:0] == 2'd2) && (bg1_color[7:0] != 8'h00)) ? bg1_color[7:0] :
           (((bg0_priority[1:0] == 2'd2) && (bg0_color[7:0] != 8'h00)) ? bg0_color[7:0] :
           (((spr_priority[1:0] == 2'd2) && (spr_color[7:0] != 8'h00)) ? spr_color[7:0] :

           // Priority 3
           (((bmp_priority[1:0] == 2'd3) && (bmp_color != 8'h00)) ? bmp_color[7:0] :
           (((bg1_priority[1:0] == 2'd3) && (bg1_color != 8'h00)) ? bg1_color[7:0] :
           (((bg0_priority[1:0] == 2'd3) && (bg0_color != 8'h00)) ? bg0_color[7:0] :
           (((spr_priority[1:0] == 2'd3) && (spr_color != 8'h00)) ? spr_color[7:0] :

           // Default to color 0 (typically black) if no layers active
           8'h00 ))))))))))))))));

    
    wire [23:0] pixel_val;
    palette_ram palram(
        .clka(cpu_clk),
        .wea(vga_pal_wea),
        .addra(cpu_addr[9:2]),
        .dina(cpu_din[23:0]),
        .clkb(!vga_clk),
        .addrb(pixel_lut[7:0]),
        .doutb(pixel_val)
    );

    
    always @(posedge vga_clk)
    begin
        vga_r <= 0;
        vga_g <= 0;
        vga_b <= 0;
        if((vga_x < h_active) && (vga_y < v_active)) begin
            vga_r <= pixel_val[23:16];
            vga_g <= pixel_val[15:8];
            vga_b <= pixel_val[7:0];
        end
        cpu_hirq <= (vga_x[10:0] >= h_active[10:0]) && (vga_y[10:0] == h_irq[10:0]);
        cpu_virq <= (vga_x[10:3] == 8'd0) && (vga_y == v_active);
    end

    vga_timing vga_timing(
      .clk(vga_clk),
      .rst(vga_rst),
      .hs(vga_hs),
      .vs(vga_vs),
      .vsi(1'b0),
      .h_front(h_front),
      .h_sync(h_sync),
      .h_back(h_back),
      .h_active(h_active),
      .v_front(v_front),
      .v_sync(v_sync),
      .v_back(v_back),
      .v_active(v_active),
      .x(vga_x),
      .y(vga_y),
      .enable(vga_blank)
    );
    
endmodule
